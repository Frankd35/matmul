`timescale 1ns / 1ps

module matmul(
    input           clk,
    input           rst,

    // matrix A & B access port
    output          mab_en,      // memory enable
    output          mab_we,      // memory write enable
    output  [ 8:0]  mab_addr,    // memory address
    input   [31:0]  mab_dout,    // memory read data
    output  [31:0]  mab_din,     // memory write data

    // matrix C access port
    output          mc_en,      // memory enable
    output          mc_we,      // memory write enable
    output  [ 7:0]  mc_addr,    // memory address
    input   [31:0]  mc_dout,    // memory read data
    output  [31:0]  mc_din,     // memory write data

    output ready
);
    reg [4:0] cnt32;
    wire clk16x, clk32x;
    assign clk16x = cnt32[3:0] == 4'd0;
    assign clk32x = cnt32 == 0;
    always @(posedge clk) begin
        if (rst) begin
			oaddr <= 0;
			out <= 0;
			finish <= 0;
            cnt32 <= 0;
        end else begin
            cnt32 <= cnt32 + 1;
        end
    end

    assign mab_en = 1;
    assign mab_we = 0;
    wire row_en;
    wire [15:0] row_shifter_en, col_shifter_en; 
    // wire [15:0] col_shifter_en; 
	wire PE_clk = out ? clk : clk32x;	// for speed up
	wire shifter_clk = out ? !clk : clk;	// for speed up
    controller ctrl(.clk(clk16x), .rst(rst), .row_en(row_en), .row_shifter_en(row_shifter_en), .col_shifter_en(col_shifter_en));
    addr_gen addr_generator(.clk(clk), .rst(rst), .row_en(row_en), .addr(mab_addr));

    /* ------------------------------------------------------------------ */
    // 输入 buffer
    // clk32x 每32周期一次 代表 col 和 row 都加载完一次向量
    wire [31:0] shifter_row_0, shifter_col_0, shifter_row_1, shifter_col_1, shifter_row_2, shifter_col_2, shifter_row_3, shifter_col_3, shifter_row_4, shifter_col_4, shifter_row_5, shifter_col_5,
    shifter_row_6, shifter_col_6, shifter_row_7, shifter_col_7, shifter_row_8, shifter_col_8, shifter_row_9, shifter_col_9, shifter_row_10, shifter_col_10, shifter_row_11, shifter_col_11, shifter_row_12,
    shifter_col_12, shifter_row_13, shifter_col_13, shifter_row_14, shifter_col_14, shifter_row_15, shifter_col_15;    

    shifter row_0(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[0]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_0));
    shifter col_0(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[0]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_0));
    shifter row_1(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[1]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_1));
    shifter col_1(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[1]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_1));
    shifter row_2(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[2]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_2));
    shifter col_2(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[2]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_2));
    shifter row_3(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[3]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_3));
    shifter col_3(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[3]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_3));
    shifter row_4(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[4]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_4));
    shifter col_4(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[4]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_4));
    shifter row_5(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[5]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_5));
    shifter col_5(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[5]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_5));
    shifter row_6(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[6]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_6));
    shifter col_6(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[6]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_6));
    shifter row_7(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[7]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_7));
    shifter col_7(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[7]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_7));
    shifter row_8(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[8]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_8));
    shifter col_8(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[8]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_8));
    shifter row_9(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[9]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_9));
    shifter col_9(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[9]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_9));
    shifter row_10(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[10]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_10));
    shifter col_10(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[10]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_10));
    shifter row_11(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[11]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_11));
    shifter col_11(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[11]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_11));
    shifter row_12(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[12]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_12));
    shifter col_12(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[12]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_12));
    shifter row_13(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[13]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_13));
    shifter col_13(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[13]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_13));
    shifter row_14(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[14]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_14));
    shifter col_14(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[14]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_14));
    shifter row_15(.clk(shifter_clk), .rst(rst), .load(row_shifter_en[15]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_row_15));
    shifter col_15(.clk(shifter_clk), .rst(rst), .load(col_shifter_en[15]), .en(out ? 1 : clk32x), .idata(mab_dout), .out(shifter_col_15));


    /* ------------------------------------------------------------------ */
    // systolic array --- 16x16 PE
	wire [31:0] sa_out [255:0];
	wire [31:0] sa_0_0_row, sa_0_0_col, 
	sa_0_1_row, sa_0_1_col, sa_0_2_row, sa_0_2_col, sa_0_3_row, sa_0_3_col, sa_0_4_row, sa_0_4_col, 
	sa_0_5_row, sa_0_5_col, sa_0_6_row, sa_0_6_col, sa_0_7_row, sa_0_7_col, sa_0_8_row, sa_0_8_col, 
	sa_0_9_row, sa_0_9_col, sa_0_10_row, sa_0_10_col, sa_0_11_row, sa_0_11_col, sa_0_12_row, sa_0_12_col, 
	sa_0_13_row, sa_0_13_col, sa_0_14_row, sa_0_14_col, sa_0_15_row, sa_0_15_col, sa_1_0_row, sa_1_0_col, 
	sa_1_1_row, sa_1_1_col, sa_1_2_row, sa_1_2_col, sa_1_3_row, sa_1_3_col, sa_1_4_row, sa_1_4_col, 
	sa_1_5_row, sa_1_5_col, sa_1_6_row, sa_1_6_col, sa_1_7_row, sa_1_7_col, sa_1_8_row, sa_1_8_col, 
	sa_1_9_row, sa_1_9_col, sa_1_10_row, sa_1_10_col, sa_1_11_row, sa_1_11_col, sa_1_12_row, sa_1_12_col, 
	sa_1_13_row, sa_1_13_col, sa_1_14_row, sa_1_14_col, sa_1_15_row, sa_1_15_col, sa_2_0_row, sa_2_0_col, 
	sa_2_1_row, sa_2_1_col, sa_2_2_row, sa_2_2_col, sa_2_3_row, sa_2_3_col, sa_2_4_row, sa_2_4_col, 
	sa_2_5_row, sa_2_5_col, sa_2_6_row, sa_2_6_col, sa_2_7_row, sa_2_7_col, sa_2_8_row, sa_2_8_col, 
	sa_2_9_row, sa_2_9_col, sa_2_10_row, sa_2_10_col, sa_2_11_row, sa_2_11_col, sa_2_12_row, sa_2_12_col, 
	sa_2_13_row, sa_2_13_col, sa_2_14_row, sa_2_14_col, sa_2_15_row, sa_2_15_col, sa_3_0_row, sa_3_0_col, 
	sa_3_1_row, sa_3_1_col, sa_3_2_row, sa_3_2_col, sa_3_3_row, sa_3_3_col, sa_3_4_row, sa_3_4_col, 
	sa_3_5_row, sa_3_5_col, sa_3_6_row, sa_3_6_col, sa_3_7_row, sa_3_7_col, sa_3_8_row, sa_3_8_col, 
	sa_3_9_row, sa_3_9_col, sa_3_10_row, sa_3_10_col, sa_3_11_row, sa_3_11_col, sa_3_12_row, sa_3_12_col, 
	sa_3_13_row, sa_3_13_col, sa_3_14_row, sa_3_14_col, sa_3_15_row, sa_3_15_col, sa_4_0_row, sa_4_0_col, 
	sa_4_1_row, sa_4_1_col, sa_4_2_row, sa_4_2_col, sa_4_3_row, sa_4_3_col, sa_4_4_row, sa_4_4_col, 
	sa_4_5_row, sa_4_5_col, sa_4_6_row, sa_4_6_col, sa_4_7_row, sa_4_7_col, sa_4_8_row, sa_4_8_col, 
	sa_4_9_row, sa_4_9_col, sa_4_10_row, sa_4_10_col, sa_4_11_row, sa_4_11_col, sa_4_12_row, sa_4_12_col, 
	sa_4_13_row, sa_4_13_col, sa_4_14_row, sa_4_14_col, sa_4_15_row, sa_4_15_col, sa_5_0_row, sa_5_0_col, 
	sa_5_1_row, sa_5_1_col, sa_5_2_row, sa_5_2_col, sa_5_3_row, sa_5_3_col, sa_5_4_row, sa_5_4_col, 
	sa_5_5_row, sa_5_5_col, sa_5_6_row, sa_5_6_col, sa_5_7_row, sa_5_7_col, sa_5_8_row, sa_5_8_col, 
	sa_5_9_row, sa_5_9_col, sa_5_10_row, sa_5_10_col, sa_5_11_row, sa_5_11_col, sa_5_12_row, sa_5_12_col, 
	sa_5_13_row, sa_5_13_col, sa_5_14_row, sa_5_14_col, sa_5_15_row, sa_5_15_col, sa_6_0_row, sa_6_0_col, 
	sa_6_1_row, sa_6_1_col, sa_6_2_row, sa_6_2_col, sa_6_3_row, sa_6_3_col, sa_6_4_row, sa_6_4_col, 
	sa_6_5_row, sa_6_5_col, sa_6_6_row, sa_6_6_col, sa_6_7_row, sa_6_7_col, sa_6_8_row, sa_6_8_col, 
	sa_6_9_row, sa_6_9_col, sa_6_10_row, sa_6_10_col, sa_6_11_row, sa_6_11_col, sa_6_12_row, sa_6_12_col, 
	sa_6_13_row, sa_6_13_col, sa_6_14_row, sa_6_14_col, sa_6_15_row, sa_6_15_col, sa_7_0_row, sa_7_0_col, 
	sa_7_1_row, sa_7_1_col, sa_7_2_row, sa_7_2_col, sa_7_3_row, sa_7_3_col, sa_7_4_row, sa_7_4_col, 
	sa_7_5_row, sa_7_5_col, sa_7_6_row, sa_7_6_col, sa_7_7_row, sa_7_7_col, sa_7_8_row, sa_7_8_col, 
	sa_7_9_row, sa_7_9_col, sa_7_10_row, sa_7_10_col, sa_7_11_row, sa_7_11_col, sa_7_12_row, sa_7_12_col, 
	sa_7_13_row, sa_7_13_col, sa_7_14_row, sa_7_14_col, sa_7_15_row, sa_7_15_col, sa_8_0_row, sa_8_0_col, 
	sa_8_1_row, sa_8_1_col, sa_8_2_row, sa_8_2_col, sa_8_3_row, sa_8_3_col, sa_8_4_row, sa_8_4_col, 
	sa_8_5_row, sa_8_5_col, sa_8_6_row, sa_8_6_col, sa_8_7_row, sa_8_7_col, sa_8_8_row, sa_8_8_col, 
	sa_8_9_row, sa_8_9_col, sa_8_10_row, sa_8_10_col, sa_8_11_row, sa_8_11_col, sa_8_12_row, sa_8_12_col, 
	sa_8_13_row, sa_8_13_col, sa_8_14_row, sa_8_14_col, sa_8_15_row, sa_8_15_col, sa_9_0_row, sa_9_0_col, 
	sa_9_1_row, sa_9_1_col, sa_9_2_row, sa_9_2_col, sa_9_3_row, sa_9_3_col, sa_9_4_row, sa_9_4_col, 
	sa_9_5_row, sa_9_5_col, sa_9_6_row, sa_9_6_col, sa_9_7_row, sa_9_7_col, sa_9_8_row, sa_9_8_col, 
	sa_9_9_row, sa_9_9_col, sa_9_10_row, sa_9_10_col, sa_9_11_row, sa_9_11_col, sa_9_12_row, sa_9_12_col, 
	sa_9_13_row, sa_9_13_col, sa_9_14_row, sa_9_14_col, sa_9_15_row, sa_9_15_col, sa_10_0_row, sa_10_0_col, 
	sa_10_1_row, sa_10_1_col, sa_10_2_row, sa_10_2_col, sa_10_3_row, sa_10_3_col, sa_10_4_row, sa_10_4_col, 
	sa_10_5_row, sa_10_5_col, sa_10_6_row, sa_10_6_col, sa_10_7_row, sa_10_7_col, sa_10_8_row, sa_10_8_col, 
	sa_10_9_row, sa_10_9_col, sa_10_10_row, sa_10_10_col, sa_10_11_row, sa_10_11_col, sa_10_12_row, sa_10_12_col, 
	sa_10_13_row, sa_10_13_col, sa_10_14_row, sa_10_14_col, sa_10_15_row, sa_10_15_col, sa_11_0_row, sa_11_0_col, 
	sa_11_1_row, sa_11_1_col, sa_11_2_row, sa_11_2_col, sa_11_3_row, sa_11_3_col, sa_11_4_row, sa_11_4_col, 
	sa_11_5_row, sa_11_5_col, sa_11_6_row, sa_11_6_col, sa_11_7_row, sa_11_7_col, sa_11_8_row, sa_11_8_col, 
	sa_11_9_row, sa_11_9_col, sa_11_10_row, sa_11_10_col, sa_11_11_row, sa_11_11_col, sa_11_12_row, sa_11_12_col, 
	sa_11_13_row, sa_11_13_col, sa_11_14_row, sa_11_14_col, sa_11_15_row, sa_11_15_col, sa_12_0_row, sa_12_0_col, 
	sa_12_1_row, sa_12_1_col, sa_12_2_row, sa_12_2_col, sa_12_3_row, sa_12_3_col, sa_12_4_row, sa_12_4_col, 
	sa_12_5_row, sa_12_5_col, sa_12_6_row, sa_12_6_col, sa_12_7_row, sa_12_7_col, sa_12_8_row, sa_12_8_col, 
	sa_12_9_row, sa_12_9_col, sa_12_10_row, sa_12_10_col, sa_12_11_row, sa_12_11_col, sa_12_12_row, sa_12_12_col, 
	sa_12_13_row, sa_12_13_col, sa_12_14_row, sa_12_14_col, sa_12_15_row, sa_12_15_col, sa_13_0_row, sa_13_0_col, 
	sa_13_1_row, sa_13_1_col, sa_13_2_row, sa_13_2_col, sa_13_3_row, sa_13_3_col, sa_13_4_row, sa_13_4_col, 
	sa_13_5_row, sa_13_5_col, sa_13_6_row, sa_13_6_col, sa_13_7_row, sa_13_7_col, sa_13_8_row, sa_13_8_col, 
	sa_13_9_row, sa_13_9_col, sa_13_10_row, sa_13_10_col, sa_13_11_row, sa_13_11_col, sa_13_12_row, sa_13_12_col, 
	sa_13_13_row, sa_13_13_col, sa_13_14_row, sa_13_14_col, sa_13_15_row, sa_13_15_col, sa_14_0_row, sa_14_0_col, 
	sa_14_1_row, sa_14_1_col, sa_14_2_row, sa_14_2_col, sa_14_3_row, sa_14_3_col, sa_14_4_row, sa_14_4_col, 
	sa_14_5_row, sa_14_5_col, sa_14_6_row, sa_14_6_col, sa_14_7_row, sa_14_7_col, sa_14_8_row, sa_14_8_col, 
	sa_14_9_row, sa_14_9_col, sa_14_10_row, sa_14_10_col, sa_14_11_row, sa_14_11_col, sa_14_12_row, sa_14_12_col, 
	sa_14_13_row, sa_14_13_col, sa_14_14_row, sa_14_14_col, sa_14_15_row, sa_14_15_col, sa_15_0_row, sa_15_0_col, 
	sa_15_1_row, sa_15_1_col, sa_15_2_row, sa_15_2_col, sa_15_3_row, sa_15_3_col, sa_15_4_row, sa_15_4_col, 
	sa_15_5_row, sa_15_5_col, sa_15_6_row, sa_15_6_col, sa_15_7_row, sa_15_7_col, sa_15_8_row, sa_15_8_col, 
	sa_15_9_row, sa_15_9_col, sa_15_10_row, sa_15_10_col, sa_15_11_row, sa_15_11_col, sa_15_12_row, sa_15_12_col, 
	sa_15_13_row, sa_15_13_col, sa_15_14_row, sa_15_14_col, sa_15_15_row, sa_15_15_col;

	PE sa_0_0(.clk(PE_clk), .rst(rst), .in_col(shifter_col_0), .in_row(shifter_row_0), .out_col(sa_0_0_col), .out_row(sa_0_0_row), .out_sum(sa_out[0]));
	PE sa_0_1(.clk(PE_clk), .rst(rst), .in_col(shifter_col_1), .in_row(sa_0_0_row), .out_col(sa_0_1_col), .out_row(sa_0_1_row), .out_sum(sa_out[1]));
	PE sa_0_2(.clk(PE_clk), .rst(rst), .in_col(shifter_col_2), .in_row(sa_0_1_row), .out_col(sa_0_2_col), .out_row(sa_0_2_row), .out_sum(sa_out[2]));
	PE sa_0_3(.clk(PE_clk), .rst(rst), .in_col(shifter_col_3), .in_row(sa_0_2_row), .out_col(sa_0_3_col), .out_row(sa_0_3_row), .out_sum(sa_out[3]));
	PE sa_0_4(.clk(PE_clk), .rst(rst), .in_col(shifter_col_4), .in_row(sa_0_3_row), .out_col(sa_0_4_col), .out_row(sa_0_4_row), .out_sum(sa_out[4]));
	PE sa_0_5(.clk(PE_clk), .rst(rst), .in_col(shifter_col_5), .in_row(sa_0_4_row), .out_col(sa_0_5_col), .out_row(sa_0_5_row), .out_sum(sa_out[5]));
	PE sa_0_6(.clk(PE_clk), .rst(rst), .in_col(shifter_col_6), .in_row(sa_0_5_row), .out_col(sa_0_6_col), .out_row(sa_0_6_row), .out_sum(sa_out[6]));
	PE sa_0_7(.clk(PE_clk), .rst(rst), .in_col(shifter_col_7), .in_row(sa_0_6_row), .out_col(sa_0_7_col), .out_row(sa_0_7_row), .out_sum(sa_out[7]));
	PE sa_0_8(.clk(PE_clk), .rst(rst), .in_col(shifter_col_8), .in_row(sa_0_7_row), .out_col(sa_0_8_col), .out_row(sa_0_8_row), .out_sum(sa_out[8]));
	PE sa_0_9(.clk(PE_clk), .rst(rst), .in_col(shifter_col_9), .in_row(sa_0_8_row), .out_col(sa_0_9_col), .out_row(sa_0_9_row), .out_sum(sa_out[9]));
	PE sa_0_10(.clk(PE_clk), .rst(rst), .in_col(shifter_col_10), .in_row(sa_0_9_row), .out_col(sa_0_10_col), .out_row(sa_0_10_row), .out_sum(sa_out[10]));
	PE sa_0_11(.clk(PE_clk), .rst(rst), .in_col(shifter_col_11), .in_row(sa_0_10_row), .out_col(sa_0_11_col), .out_row(sa_0_11_row), .out_sum(sa_out[11]));
	PE sa_0_12(.clk(PE_clk), .rst(rst), .in_col(shifter_col_12), .in_row(sa_0_11_row), .out_col(sa_0_12_col), .out_row(sa_0_12_row), .out_sum(sa_out[12]));
	PE sa_0_13(.clk(PE_clk), .rst(rst), .in_col(shifter_col_13), .in_row(sa_0_12_row), .out_col(sa_0_13_col), .out_row(sa_0_13_row), .out_sum(sa_out[13]));
	PE sa_0_14(.clk(PE_clk), .rst(rst), .in_col(shifter_col_14), .in_row(sa_0_13_row), .out_col(sa_0_14_col), .out_row(sa_0_14_row), .out_sum(sa_out[14]));
	PE sa_0_15(.clk(PE_clk), .rst(rst), .in_col(shifter_col_15), .in_row(sa_0_14_row), .out_col(sa_0_15_col), .out_row(sa_0_15_row), .out_sum(sa_out[15]));
	PE sa_1_0(.clk(PE_clk), .rst(rst), .in_col(sa_0_0_col), .in_row(shifter_row_1), .out_col(sa_1_0_col), .out_row(sa_1_0_row), .out_sum(sa_out[16]));
	PE sa_1_1(.clk(PE_clk), .rst(rst), .in_col(sa_0_1_col), .in_row(sa_1_0_row), .out_col(sa_1_1_col), .out_row(sa_1_1_row), .out_sum(sa_out[17]));
	PE sa_1_2(.clk(PE_clk), .rst(rst), .in_col(sa_0_2_col), .in_row(sa_1_1_row), .out_col(sa_1_2_col), .out_row(sa_1_2_row), .out_sum(sa_out[18]));
	PE sa_1_3(.clk(PE_clk), .rst(rst), .in_col(sa_0_3_col), .in_row(sa_1_2_row), .out_col(sa_1_3_col), .out_row(sa_1_3_row), .out_sum(sa_out[19]));
	PE sa_1_4(.clk(PE_clk), .rst(rst), .in_col(sa_0_4_col), .in_row(sa_1_3_row), .out_col(sa_1_4_col), .out_row(sa_1_4_row), .out_sum(sa_out[20]));
	PE sa_1_5(.clk(PE_clk), .rst(rst), .in_col(sa_0_5_col), .in_row(sa_1_4_row), .out_col(sa_1_5_col), .out_row(sa_1_5_row), .out_sum(sa_out[21]));
	PE sa_1_6(.clk(PE_clk), .rst(rst), .in_col(sa_0_6_col), .in_row(sa_1_5_row), .out_col(sa_1_6_col), .out_row(sa_1_6_row), .out_sum(sa_out[22]));
	PE sa_1_7(.clk(PE_clk), .rst(rst), .in_col(sa_0_7_col), .in_row(sa_1_6_row), .out_col(sa_1_7_col), .out_row(sa_1_7_row), .out_sum(sa_out[23]));
	PE sa_1_8(.clk(PE_clk), .rst(rst), .in_col(sa_0_8_col), .in_row(sa_1_7_row), .out_col(sa_1_8_col), .out_row(sa_1_8_row), .out_sum(sa_out[24]));
	PE sa_1_9(.clk(PE_clk), .rst(rst), .in_col(sa_0_9_col), .in_row(sa_1_8_row), .out_col(sa_1_9_col), .out_row(sa_1_9_row), .out_sum(sa_out[25]));
	PE sa_1_10(.clk(PE_clk), .rst(rst), .in_col(sa_0_10_col), .in_row(sa_1_9_row), .out_col(sa_1_10_col), .out_row(sa_1_10_row), .out_sum(sa_out[26]));
	PE sa_1_11(.clk(PE_clk), .rst(rst), .in_col(sa_0_11_col), .in_row(sa_1_10_row), .out_col(sa_1_11_col), .out_row(sa_1_11_row), .out_sum(sa_out[27]));
	PE sa_1_12(.clk(PE_clk), .rst(rst), .in_col(sa_0_12_col), .in_row(sa_1_11_row), .out_col(sa_1_12_col), .out_row(sa_1_12_row), .out_sum(sa_out[28]));
	PE sa_1_13(.clk(PE_clk), .rst(rst), .in_col(sa_0_13_col), .in_row(sa_1_12_row), .out_col(sa_1_13_col), .out_row(sa_1_13_row), .out_sum(sa_out[29]));
	PE sa_1_14(.clk(PE_clk), .rst(rst), .in_col(sa_0_14_col), .in_row(sa_1_13_row), .out_col(sa_1_14_col), .out_row(sa_1_14_row), .out_sum(sa_out[30]));
	PE sa_1_15(.clk(PE_clk), .rst(rst), .in_col(sa_0_15_col), .in_row(sa_1_14_row), .out_col(sa_1_15_col), .out_row(sa_1_15_row), .out_sum(sa_out[31]));
	PE sa_2_0(.clk(PE_clk), .rst(rst), .in_col(sa_1_0_col), .in_row(shifter_row_2), .out_col(sa_2_0_col), .out_row(sa_2_0_row), .out_sum(sa_out[32]));
	PE sa_2_1(.clk(PE_clk), .rst(rst), .in_col(sa_1_1_col), .in_row(sa_2_0_row), .out_col(sa_2_1_col), .out_row(sa_2_1_row), .out_sum(sa_out[33]));
	PE sa_2_2(.clk(PE_clk), .rst(rst), .in_col(sa_1_2_col), .in_row(sa_2_1_row), .out_col(sa_2_2_col), .out_row(sa_2_2_row), .out_sum(sa_out[34]));
	PE sa_2_3(.clk(PE_clk), .rst(rst), .in_col(sa_1_3_col), .in_row(sa_2_2_row), .out_col(sa_2_3_col), .out_row(sa_2_3_row), .out_sum(sa_out[35]));
	PE sa_2_4(.clk(PE_clk), .rst(rst), .in_col(sa_1_4_col), .in_row(sa_2_3_row), .out_col(sa_2_4_col), .out_row(sa_2_4_row), .out_sum(sa_out[36]));
	PE sa_2_5(.clk(PE_clk), .rst(rst), .in_col(sa_1_5_col), .in_row(sa_2_4_row), .out_col(sa_2_5_col), .out_row(sa_2_5_row), .out_sum(sa_out[37]));
	PE sa_2_6(.clk(PE_clk), .rst(rst), .in_col(sa_1_6_col), .in_row(sa_2_5_row), .out_col(sa_2_6_col), .out_row(sa_2_6_row), .out_sum(sa_out[38]));
	PE sa_2_7(.clk(PE_clk), .rst(rst), .in_col(sa_1_7_col), .in_row(sa_2_6_row), .out_col(sa_2_7_col), .out_row(sa_2_7_row), .out_sum(sa_out[39]));
	PE sa_2_8(.clk(PE_clk), .rst(rst), .in_col(sa_1_8_col), .in_row(sa_2_7_row), .out_col(sa_2_8_col), .out_row(sa_2_8_row), .out_sum(sa_out[40]));
	PE sa_2_9(.clk(PE_clk), .rst(rst), .in_col(sa_1_9_col), .in_row(sa_2_8_row), .out_col(sa_2_9_col), .out_row(sa_2_9_row), .out_sum(sa_out[41]));
	PE sa_2_10(.clk(PE_clk), .rst(rst), .in_col(sa_1_10_col), .in_row(sa_2_9_row), .out_col(sa_2_10_col), .out_row(sa_2_10_row), .out_sum(sa_out[42]));
	PE sa_2_11(.clk(PE_clk), .rst(rst), .in_col(sa_1_11_col), .in_row(sa_2_10_row), .out_col(sa_2_11_col), .out_row(sa_2_11_row), .out_sum(sa_out[43]));
	PE sa_2_12(.clk(PE_clk), .rst(rst), .in_col(sa_1_12_col), .in_row(sa_2_11_row), .out_col(sa_2_12_col), .out_row(sa_2_12_row), .out_sum(sa_out[44]));
	PE sa_2_13(.clk(PE_clk), .rst(rst), .in_col(sa_1_13_col), .in_row(sa_2_12_row), .out_col(sa_2_13_col), .out_row(sa_2_13_row), .out_sum(sa_out[45]));
	PE sa_2_14(.clk(PE_clk), .rst(rst), .in_col(sa_1_14_col), .in_row(sa_2_13_row), .out_col(sa_2_14_col), .out_row(sa_2_14_row), .out_sum(sa_out[46]));
	PE sa_2_15(.clk(PE_clk), .rst(rst), .in_col(sa_1_15_col), .in_row(sa_2_14_row), .out_col(sa_2_15_col), .out_row(sa_2_15_row), .out_sum(sa_out[47]));
	PE sa_3_0(.clk(PE_clk), .rst(rst), .in_col(sa_2_0_col), .in_row(shifter_row_3), .out_col(sa_3_0_col), .out_row(sa_3_0_row), .out_sum(sa_out[48]));
	PE sa_3_1(.clk(PE_clk), .rst(rst), .in_col(sa_2_1_col), .in_row(sa_3_0_row), .out_col(sa_3_1_col), .out_row(sa_3_1_row), .out_sum(sa_out[49]));
	PE sa_3_2(.clk(PE_clk), .rst(rst), .in_col(sa_2_2_col), .in_row(sa_3_1_row), .out_col(sa_3_2_col), .out_row(sa_3_2_row), .out_sum(sa_out[50]));
	PE sa_3_3(.clk(PE_clk), .rst(rst), .in_col(sa_2_3_col), .in_row(sa_3_2_row), .out_col(sa_3_3_col), .out_row(sa_3_3_row), .out_sum(sa_out[51]));
	PE sa_3_4(.clk(PE_clk), .rst(rst), .in_col(sa_2_4_col), .in_row(sa_3_3_row), .out_col(sa_3_4_col), .out_row(sa_3_4_row), .out_sum(sa_out[52]));
	PE sa_3_5(.clk(PE_clk), .rst(rst), .in_col(sa_2_5_col), .in_row(sa_3_4_row), .out_col(sa_3_5_col), .out_row(sa_3_5_row), .out_sum(sa_out[53]));
	PE sa_3_6(.clk(PE_clk), .rst(rst), .in_col(sa_2_6_col), .in_row(sa_3_5_row), .out_col(sa_3_6_col), .out_row(sa_3_6_row), .out_sum(sa_out[54]));
	PE sa_3_7(.clk(PE_clk), .rst(rst), .in_col(sa_2_7_col), .in_row(sa_3_6_row), .out_col(sa_3_7_col), .out_row(sa_3_7_row), .out_sum(sa_out[55]));
	PE sa_3_8(.clk(PE_clk), .rst(rst), .in_col(sa_2_8_col), .in_row(sa_3_7_row), .out_col(sa_3_8_col), .out_row(sa_3_8_row), .out_sum(sa_out[56]));
	PE sa_3_9(.clk(PE_clk), .rst(rst), .in_col(sa_2_9_col), .in_row(sa_3_8_row), .out_col(sa_3_9_col), .out_row(sa_3_9_row), .out_sum(sa_out[57]));
	PE sa_3_10(.clk(PE_clk), .rst(rst), .in_col(sa_2_10_col), .in_row(sa_3_9_row), .out_col(sa_3_10_col), .out_row(sa_3_10_row), .out_sum(sa_out[58]));
	PE sa_3_11(.clk(PE_clk), .rst(rst), .in_col(sa_2_11_col), .in_row(sa_3_10_row), .out_col(sa_3_11_col), .out_row(sa_3_11_row), .out_sum(sa_out[59]));
	PE sa_3_12(.clk(PE_clk), .rst(rst), .in_col(sa_2_12_col), .in_row(sa_3_11_row), .out_col(sa_3_12_col), .out_row(sa_3_12_row), .out_sum(sa_out[60]));
	PE sa_3_13(.clk(PE_clk), .rst(rst), .in_col(sa_2_13_col), .in_row(sa_3_12_row), .out_col(sa_3_13_col), .out_row(sa_3_13_row), .out_sum(sa_out[61]));
	PE sa_3_14(.clk(PE_clk), .rst(rst), .in_col(sa_2_14_col), .in_row(sa_3_13_row), .out_col(sa_3_14_col), .out_row(sa_3_14_row), .out_sum(sa_out[62]));
	PE sa_3_15(.clk(PE_clk), .rst(rst), .in_col(sa_2_15_col), .in_row(sa_3_14_row), .out_col(sa_3_15_col), .out_row(sa_3_15_row), .out_sum(sa_out[63]));
	PE sa_4_0(.clk(PE_clk), .rst(rst), .in_col(sa_3_0_col), .in_row(shifter_row_4), .out_col(sa_4_0_col), .out_row(sa_4_0_row), .out_sum(sa_out[64]));
	PE sa_4_1(.clk(PE_clk), .rst(rst), .in_col(sa_3_1_col), .in_row(sa_4_0_row), .out_col(sa_4_1_col), .out_row(sa_4_1_row), .out_sum(sa_out[65]));
	PE sa_4_2(.clk(PE_clk), .rst(rst), .in_col(sa_3_2_col), .in_row(sa_4_1_row), .out_col(sa_4_2_col), .out_row(sa_4_2_row), .out_sum(sa_out[66]));
	PE sa_4_3(.clk(PE_clk), .rst(rst), .in_col(sa_3_3_col), .in_row(sa_4_2_row), .out_col(sa_4_3_col), .out_row(sa_4_3_row), .out_sum(sa_out[67]));
	PE sa_4_4(.clk(PE_clk), .rst(rst), .in_col(sa_3_4_col), .in_row(sa_4_3_row), .out_col(sa_4_4_col), .out_row(sa_4_4_row), .out_sum(sa_out[68]));
	PE sa_4_5(.clk(PE_clk), .rst(rst), .in_col(sa_3_5_col), .in_row(sa_4_4_row), .out_col(sa_4_5_col), .out_row(sa_4_5_row), .out_sum(sa_out[69]));
	PE sa_4_6(.clk(PE_clk), .rst(rst), .in_col(sa_3_6_col), .in_row(sa_4_5_row), .out_col(sa_4_6_col), .out_row(sa_4_6_row), .out_sum(sa_out[70]));
	PE sa_4_7(.clk(PE_clk), .rst(rst), .in_col(sa_3_7_col), .in_row(sa_4_6_row), .out_col(sa_4_7_col), .out_row(sa_4_7_row), .out_sum(sa_out[71]));
	PE sa_4_8(.clk(PE_clk), .rst(rst), .in_col(sa_3_8_col), .in_row(sa_4_7_row), .out_col(sa_4_8_col), .out_row(sa_4_8_row), .out_sum(sa_out[72]));
	PE sa_4_9(.clk(PE_clk), .rst(rst), .in_col(sa_3_9_col), .in_row(sa_4_8_row), .out_col(sa_4_9_col), .out_row(sa_4_9_row), .out_sum(sa_out[73]));
	PE sa_4_10(.clk(PE_clk), .rst(rst), .in_col(sa_3_10_col), .in_row(sa_4_9_row), .out_col(sa_4_10_col), .out_row(sa_4_10_row), .out_sum(sa_out[74]));
	PE sa_4_11(.clk(PE_clk), .rst(rst), .in_col(sa_3_11_col), .in_row(sa_4_10_row), .out_col(sa_4_11_col), .out_row(sa_4_11_row), .out_sum(sa_out[75]));
	PE sa_4_12(.clk(PE_clk), .rst(rst), .in_col(sa_3_12_col), .in_row(sa_4_11_row), .out_col(sa_4_12_col), .out_row(sa_4_12_row), .out_sum(sa_out[76]));
	PE sa_4_13(.clk(PE_clk), .rst(rst), .in_col(sa_3_13_col), .in_row(sa_4_12_row), .out_col(sa_4_13_col), .out_row(sa_4_13_row), .out_sum(sa_out[77]));
	PE sa_4_14(.clk(PE_clk), .rst(rst), .in_col(sa_3_14_col), .in_row(sa_4_13_row), .out_col(sa_4_14_col), .out_row(sa_4_14_row), .out_sum(sa_out[78]));
	PE sa_4_15(.clk(PE_clk), .rst(rst), .in_col(sa_3_15_col), .in_row(sa_4_14_row), .out_col(sa_4_15_col), .out_row(sa_4_15_row), .out_sum(sa_out[79]));
	PE sa_5_0(.clk(PE_clk), .rst(rst), .in_col(sa_4_0_col), .in_row(shifter_row_5), .out_col(sa_5_0_col), .out_row(sa_5_0_row), .out_sum(sa_out[80]));
	PE sa_5_1(.clk(PE_clk), .rst(rst), .in_col(sa_4_1_col), .in_row(sa_5_0_row), .out_col(sa_5_1_col), .out_row(sa_5_1_row), .out_sum(sa_out[81]));
	PE sa_5_2(.clk(PE_clk), .rst(rst), .in_col(sa_4_2_col), .in_row(sa_5_1_row), .out_col(sa_5_2_col), .out_row(sa_5_2_row), .out_sum(sa_out[82]));
	PE sa_5_3(.clk(PE_clk), .rst(rst), .in_col(sa_4_3_col), .in_row(sa_5_2_row), .out_col(sa_5_3_col), .out_row(sa_5_3_row), .out_sum(sa_out[83]));
	PE sa_5_4(.clk(PE_clk), .rst(rst), .in_col(sa_4_4_col), .in_row(sa_5_3_row), .out_col(sa_5_4_col), .out_row(sa_5_4_row), .out_sum(sa_out[84]));
	PE sa_5_5(.clk(PE_clk), .rst(rst), .in_col(sa_4_5_col), .in_row(sa_5_4_row), .out_col(sa_5_5_col), .out_row(sa_5_5_row), .out_sum(sa_out[85]));
	PE sa_5_6(.clk(PE_clk), .rst(rst), .in_col(sa_4_6_col), .in_row(sa_5_5_row), .out_col(sa_5_6_col), .out_row(sa_5_6_row), .out_sum(sa_out[86]));
	PE sa_5_7(.clk(PE_clk), .rst(rst), .in_col(sa_4_7_col), .in_row(sa_5_6_row), .out_col(sa_5_7_col), .out_row(sa_5_7_row), .out_sum(sa_out[87]));
	PE sa_5_8(.clk(PE_clk), .rst(rst), .in_col(sa_4_8_col), .in_row(sa_5_7_row), .out_col(sa_5_8_col), .out_row(sa_5_8_row), .out_sum(sa_out[88]));
	PE sa_5_9(.clk(PE_clk), .rst(rst), .in_col(sa_4_9_col), .in_row(sa_5_8_row), .out_col(sa_5_9_col), .out_row(sa_5_9_row), .out_sum(sa_out[89]));
	PE sa_5_10(.clk(PE_clk), .rst(rst), .in_col(sa_4_10_col), .in_row(sa_5_9_row), .out_col(sa_5_10_col), .out_row(sa_5_10_row), .out_sum(sa_out[90]));
	PE sa_5_11(.clk(PE_clk), .rst(rst), .in_col(sa_4_11_col), .in_row(sa_5_10_row), .out_col(sa_5_11_col), .out_row(sa_5_11_row), .out_sum(sa_out[91]));
	PE sa_5_12(.clk(PE_clk), .rst(rst), .in_col(sa_4_12_col), .in_row(sa_5_11_row), .out_col(sa_5_12_col), .out_row(sa_5_12_row), .out_sum(sa_out[92]));
	PE sa_5_13(.clk(PE_clk), .rst(rst), .in_col(sa_4_13_col), .in_row(sa_5_12_row), .out_col(sa_5_13_col), .out_row(sa_5_13_row), .out_sum(sa_out[93]));
	PE sa_5_14(.clk(PE_clk), .rst(rst), .in_col(sa_4_14_col), .in_row(sa_5_13_row), .out_col(sa_5_14_col), .out_row(sa_5_14_row), .out_sum(sa_out[94]));
	PE sa_5_15(.clk(PE_clk), .rst(rst), .in_col(sa_4_15_col), .in_row(sa_5_14_row), .out_col(sa_5_15_col), .out_row(sa_5_15_row), .out_sum(sa_out[95]));
	PE sa_6_0(.clk(PE_clk), .rst(rst), .in_col(sa_5_0_col), .in_row(shifter_row_6), .out_col(sa_6_0_col), .out_row(sa_6_0_row), .out_sum(sa_out[96]));
	PE sa_6_1(.clk(PE_clk), .rst(rst), .in_col(sa_5_1_col), .in_row(sa_6_0_row), .out_col(sa_6_1_col), .out_row(sa_6_1_row), .out_sum(sa_out[97]));
	PE sa_6_2(.clk(PE_clk), .rst(rst), .in_col(sa_5_2_col), .in_row(sa_6_1_row), .out_col(sa_6_2_col), .out_row(sa_6_2_row), .out_sum(sa_out[98]));
	PE sa_6_3(.clk(PE_clk), .rst(rst), .in_col(sa_5_3_col), .in_row(sa_6_2_row), .out_col(sa_6_3_col), .out_row(sa_6_3_row), .out_sum(sa_out[99]));
	PE sa_6_4(.clk(PE_clk), .rst(rst), .in_col(sa_5_4_col), .in_row(sa_6_3_row), .out_col(sa_6_4_col), .out_row(sa_6_4_row), .out_sum(sa_out[100]));
	PE sa_6_5(.clk(PE_clk), .rst(rst), .in_col(sa_5_5_col), .in_row(sa_6_4_row), .out_col(sa_6_5_col), .out_row(sa_6_5_row), .out_sum(sa_out[101]));
	PE sa_6_6(.clk(PE_clk), .rst(rst), .in_col(sa_5_6_col), .in_row(sa_6_5_row), .out_col(sa_6_6_col), .out_row(sa_6_6_row), .out_sum(sa_out[102]));
	PE sa_6_7(.clk(PE_clk), .rst(rst), .in_col(sa_5_7_col), .in_row(sa_6_6_row), .out_col(sa_6_7_col), .out_row(sa_6_7_row), .out_sum(sa_out[103]));
	PE sa_6_8(.clk(PE_clk), .rst(rst), .in_col(sa_5_8_col), .in_row(sa_6_7_row), .out_col(sa_6_8_col), .out_row(sa_6_8_row), .out_sum(sa_out[104]));
	PE sa_6_9(.clk(PE_clk), .rst(rst), .in_col(sa_5_9_col), .in_row(sa_6_8_row), .out_col(sa_6_9_col), .out_row(sa_6_9_row), .out_sum(sa_out[105]));
	PE sa_6_10(.clk(PE_clk), .rst(rst), .in_col(sa_5_10_col), .in_row(sa_6_9_row), .out_col(sa_6_10_col), .out_row(sa_6_10_row), .out_sum(sa_out[106]));
	PE sa_6_11(.clk(PE_clk), .rst(rst), .in_col(sa_5_11_col), .in_row(sa_6_10_row), .out_col(sa_6_11_col), .out_row(sa_6_11_row), .out_sum(sa_out[107]));
	PE sa_6_12(.clk(PE_clk), .rst(rst), .in_col(sa_5_12_col), .in_row(sa_6_11_row), .out_col(sa_6_12_col), .out_row(sa_6_12_row), .out_sum(sa_out[108]));
	PE sa_6_13(.clk(PE_clk), .rst(rst), .in_col(sa_5_13_col), .in_row(sa_6_12_row), .out_col(sa_6_13_col), .out_row(sa_6_13_row), .out_sum(sa_out[109]));
	PE sa_6_14(.clk(PE_clk), .rst(rst), .in_col(sa_5_14_col), .in_row(sa_6_13_row), .out_col(sa_6_14_col), .out_row(sa_6_14_row), .out_sum(sa_out[110]));
	PE sa_6_15(.clk(PE_clk), .rst(rst), .in_col(sa_5_15_col), .in_row(sa_6_14_row), .out_col(sa_6_15_col), .out_row(sa_6_15_row), .out_sum(sa_out[111]));
	PE sa_7_0(.clk(PE_clk), .rst(rst), .in_col(sa_6_0_col), .in_row(shifter_row_7), .out_col(sa_7_0_col), .out_row(sa_7_0_row), .out_sum(sa_out[112]));
	PE sa_7_1(.clk(PE_clk), .rst(rst), .in_col(sa_6_1_col), .in_row(sa_7_0_row), .out_col(sa_7_1_col), .out_row(sa_7_1_row), .out_sum(sa_out[113]));
	PE sa_7_2(.clk(PE_clk), .rst(rst), .in_col(sa_6_2_col), .in_row(sa_7_1_row), .out_col(sa_7_2_col), .out_row(sa_7_2_row), .out_sum(sa_out[114]));
	PE sa_7_3(.clk(PE_clk), .rst(rst), .in_col(sa_6_3_col), .in_row(sa_7_2_row), .out_col(sa_7_3_col), .out_row(sa_7_3_row), .out_sum(sa_out[115]));
	PE sa_7_4(.clk(PE_clk), .rst(rst), .in_col(sa_6_4_col), .in_row(sa_7_3_row), .out_col(sa_7_4_col), .out_row(sa_7_4_row), .out_sum(sa_out[116]));
	PE sa_7_5(.clk(PE_clk), .rst(rst), .in_col(sa_6_5_col), .in_row(sa_7_4_row), .out_col(sa_7_5_col), .out_row(sa_7_5_row), .out_sum(sa_out[117]));
	PE sa_7_6(.clk(PE_clk), .rst(rst), .in_col(sa_6_6_col), .in_row(sa_7_5_row), .out_col(sa_7_6_col), .out_row(sa_7_6_row), .out_sum(sa_out[118]));
	PE sa_7_7(.clk(PE_clk), .rst(rst), .in_col(sa_6_7_col), .in_row(sa_7_6_row), .out_col(sa_7_7_col), .out_row(sa_7_7_row), .out_sum(sa_out[119]));
	PE sa_7_8(.clk(PE_clk), .rst(rst), .in_col(sa_6_8_col), .in_row(sa_7_7_row), .out_col(sa_7_8_col), .out_row(sa_7_8_row), .out_sum(sa_out[120]));
	PE sa_7_9(.clk(PE_clk), .rst(rst), .in_col(sa_6_9_col), .in_row(sa_7_8_row), .out_col(sa_7_9_col), .out_row(sa_7_9_row), .out_sum(sa_out[121]));
	PE sa_7_10(.clk(PE_clk), .rst(rst), .in_col(sa_6_10_col), .in_row(sa_7_9_row), .out_col(sa_7_10_col), .out_row(sa_7_10_row), .out_sum(sa_out[122]));
	PE sa_7_11(.clk(PE_clk), .rst(rst), .in_col(sa_6_11_col), .in_row(sa_7_10_row), .out_col(sa_7_11_col), .out_row(sa_7_11_row), .out_sum(sa_out[123]));
	PE sa_7_12(.clk(PE_clk), .rst(rst), .in_col(sa_6_12_col), .in_row(sa_7_11_row), .out_col(sa_7_12_col), .out_row(sa_7_12_row), .out_sum(sa_out[124]));
	PE sa_7_13(.clk(PE_clk), .rst(rst), .in_col(sa_6_13_col), .in_row(sa_7_12_row), .out_col(sa_7_13_col), .out_row(sa_7_13_row), .out_sum(sa_out[125]));
	PE sa_7_14(.clk(PE_clk), .rst(rst), .in_col(sa_6_14_col), .in_row(sa_7_13_row), .out_col(sa_7_14_col), .out_row(sa_7_14_row), .out_sum(sa_out[126]));
	PE sa_7_15(.clk(PE_clk), .rst(rst), .in_col(sa_6_15_col), .in_row(sa_7_14_row), .out_col(sa_7_15_col), .out_row(sa_7_15_row), .out_sum(sa_out[127]));
	PE sa_8_0(.clk(PE_clk), .rst(rst), .in_col(sa_7_0_col), .in_row(shifter_row_8), .out_col(sa_8_0_col), .out_row(sa_8_0_row), .out_sum(sa_out[128]));
	PE sa_8_1(.clk(PE_clk), .rst(rst), .in_col(sa_7_1_col), .in_row(sa_8_0_row), .out_col(sa_8_1_col), .out_row(sa_8_1_row), .out_sum(sa_out[129]));
	PE sa_8_2(.clk(PE_clk), .rst(rst), .in_col(sa_7_2_col), .in_row(sa_8_1_row), .out_col(sa_8_2_col), .out_row(sa_8_2_row), .out_sum(sa_out[130]));
	PE sa_8_3(.clk(PE_clk), .rst(rst), .in_col(sa_7_3_col), .in_row(sa_8_2_row), .out_col(sa_8_3_col), .out_row(sa_8_3_row), .out_sum(sa_out[131]));
	PE sa_8_4(.clk(PE_clk), .rst(rst), .in_col(sa_7_4_col), .in_row(sa_8_3_row), .out_col(sa_8_4_col), .out_row(sa_8_4_row), .out_sum(sa_out[132]));
	PE sa_8_5(.clk(PE_clk), .rst(rst), .in_col(sa_7_5_col), .in_row(sa_8_4_row), .out_col(sa_8_5_col), .out_row(sa_8_5_row), .out_sum(sa_out[133]));
	PE sa_8_6(.clk(PE_clk), .rst(rst), .in_col(sa_7_6_col), .in_row(sa_8_5_row), .out_col(sa_8_6_col), .out_row(sa_8_6_row), .out_sum(sa_out[134]));
	PE sa_8_7(.clk(PE_clk), .rst(rst), .in_col(sa_7_7_col), .in_row(sa_8_6_row), .out_col(sa_8_7_col), .out_row(sa_8_7_row), .out_sum(sa_out[135]));
	PE sa_8_8(.clk(PE_clk), .rst(rst), .in_col(sa_7_8_col), .in_row(sa_8_7_row), .out_col(sa_8_8_col), .out_row(sa_8_8_row), .out_sum(sa_out[136]));
	PE sa_8_9(.clk(PE_clk), .rst(rst), .in_col(sa_7_9_col), .in_row(sa_8_8_row), .out_col(sa_8_9_col), .out_row(sa_8_9_row), .out_sum(sa_out[137]));
	PE sa_8_10(.clk(PE_clk), .rst(rst), .in_col(sa_7_10_col), .in_row(sa_8_9_row), .out_col(sa_8_10_col), .out_row(sa_8_10_row), .out_sum(sa_out[138]));
	PE sa_8_11(.clk(PE_clk), .rst(rst), .in_col(sa_7_11_col), .in_row(sa_8_10_row), .out_col(sa_8_11_col), .out_row(sa_8_11_row), .out_sum(sa_out[139]));
	PE sa_8_12(.clk(PE_clk), .rst(rst), .in_col(sa_7_12_col), .in_row(sa_8_11_row), .out_col(sa_8_12_col), .out_row(sa_8_12_row), .out_sum(sa_out[140]));
	PE sa_8_13(.clk(PE_clk), .rst(rst), .in_col(sa_7_13_col), .in_row(sa_8_12_row), .out_col(sa_8_13_col), .out_row(sa_8_13_row), .out_sum(sa_out[141]));
	PE sa_8_14(.clk(PE_clk), .rst(rst), .in_col(sa_7_14_col), .in_row(sa_8_13_row), .out_col(sa_8_14_col), .out_row(sa_8_14_row), .out_sum(sa_out[142]));
	PE sa_8_15(.clk(PE_clk), .rst(rst), .in_col(sa_7_15_col), .in_row(sa_8_14_row), .out_col(sa_8_15_col), .out_row(sa_8_15_row), .out_sum(sa_out[143]));
	PE sa_9_0(.clk(PE_clk), .rst(rst), .in_col(sa_8_0_col), .in_row(shifter_row_9), .out_col(sa_9_0_col), .out_row(sa_9_0_row), .out_sum(sa_out[144]));
	PE sa_9_1(.clk(PE_clk), .rst(rst), .in_col(sa_8_1_col), .in_row(sa_9_0_row), .out_col(sa_9_1_col), .out_row(sa_9_1_row), .out_sum(sa_out[145]));
	PE sa_9_2(.clk(PE_clk), .rst(rst), .in_col(sa_8_2_col), .in_row(sa_9_1_row), .out_col(sa_9_2_col), .out_row(sa_9_2_row), .out_sum(sa_out[146]));
	PE sa_9_3(.clk(PE_clk), .rst(rst), .in_col(sa_8_3_col), .in_row(sa_9_2_row), .out_col(sa_9_3_col), .out_row(sa_9_3_row), .out_sum(sa_out[147]));
	PE sa_9_4(.clk(PE_clk), .rst(rst), .in_col(sa_8_4_col), .in_row(sa_9_3_row), .out_col(sa_9_4_col), .out_row(sa_9_4_row), .out_sum(sa_out[148]));
	PE sa_9_5(.clk(PE_clk), .rst(rst), .in_col(sa_8_5_col), .in_row(sa_9_4_row), .out_col(sa_9_5_col), .out_row(sa_9_5_row), .out_sum(sa_out[149]));
	PE sa_9_6(.clk(PE_clk), .rst(rst), .in_col(sa_8_6_col), .in_row(sa_9_5_row), .out_col(sa_9_6_col), .out_row(sa_9_6_row), .out_sum(sa_out[150]));
	PE sa_9_7(.clk(PE_clk), .rst(rst), .in_col(sa_8_7_col), .in_row(sa_9_6_row), .out_col(sa_9_7_col), .out_row(sa_9_7_row), .out_sum(sa_out[151]));
	PE sa_9_8(.clk(PE_clk), .rst(rst), .in_col(sa_8_8_col), .in_row(sa_9_7_row), .out_col(sa_9_8_col), .out_row(sa_9_8_row), .out_sum(sa_out[152]));
	PE sa_9_9(.clk(PE_clk), .rst(rst), .in_col(sa_8_9_col), .in_row(sa_9_8_row), .out_col(sa_9_9_col), .out_row(sa_9_9_row), .out_sum(sa_out[153]));
	PE sa_9_10(.clk(PE_clk), .rst(rst), .in_col(sa_8_10_col), .in_row(sa_9_9_row), .out_col(sa_9_10_col), .out_row(sa_9_10_row), .out_sum(sa_out[154]));
	PE sa_9_11(.clk(PE_clk), .rst(rst), .in_col(sa_8_11_col), .in_row(sa_9_10_row), .out_col(sa_9_11_col), .out_row(sa_9_11_row), .out_sum(sa_out[155]));
	PE sa_9_12(.clk(PE_clk), .rst(rst), .in_col(sa_8_12_col), .in_row(sa_9_11_row), .out_col(sa_9_12_col), .out_row(sa_9_12_row), .out_sum(sa_out[156]));
	PE sa_9_13(.clk(PE_clk), .rst(rst), .in_col(sa_8_13_col), .in_row(sa_9_12_row), .out_col(sa_9_13_col), .out_row(sa_9_13_row), .out_sum(sa_out[157]));
	PE sa_9_14(.clk(PE_clk), .rst(rst), .in_col(sa_8_14_col), .in_row(sa_9_13_row), .out_col(sa_9_14_col), .out_row(sa_9_14_row), .out_sum(sa_out[158]));
	PE sa_9_15(.clk(PE_clk), .rst(rst), .in_col(sa_8_15_col), .in_row(sa_9_14_row), .out_col(sa_9_15_col), .out_row(sa_9_15_row), .out_sum(sa_out[159]));
	PE sa_10_0(.clk(PE_clk), .rst(rst), .in_col(sa_9_0_col), .in_row(shifter_row_10), .out_col(sa_10_0_col), .out_row(sa_10_0_row), .out_sum(sa_out[160]));
	PE sa_10_1(.clk(PE_clk), .rst(rst), .in_col(sa_9_1_col), .in_row(sa_10_0_row), .out_col(sa_10_1_col), .out_row(sa_10_1_row), .out_sum(sa_out[161]));
	PE sa_10_2(.clk(PE_clk), .rst(rst), .in_col(sa_9_2_col), .in_row(sa_10_1_row), .out_col(sa_10_2_col), .out_row(sa_10_2_row), .out_sum(sa_out[162]));
	PE sa_10_3(.clk(PE_clk), .rst(rst), .in_col(sa_9_3_col), .in_row(sa_10_2_row), .out_col(sa_10_3_col), .out_row(sa_10_3_row), .out_sum(sa_out[163]));
	PE sa_10_4(.clk(PE_clk), .rst(rst), .in_col(sa_9_4_col), .in_row(sa_10_3_row), .out_col(sa_10_4_col), .out_row(sa_10_4_row), .out_sum(sa_out[164]));
	PE sa_10_5(.clk(PE_clk), .rst(rst), .in_col(sa_9_5_col), .in_row(sa_10_4_row), .out_col(sa_10_5_col), .out_row(sa_10_5_row), .out_sum(sa_out[165]));
	PE sa_10_6(.clk(PE_clk), .rst(rst), .in_col(sa_9_6_col), .in_row(sa_10_5_row), .out_col(sa_10_6_col), .out_row(sa_10_6_row), .out_sum(sa_out[166]));
	PE sa_10_7(.clk(PE_clk), .rst(rst), .in_col(sa_9_7_col), .in_row(sa_10_6_row), .out_col(sa_10_7_col), .out_row(sa_10_7_row), .out_sum(sa_out[167]));
	PE sa_10_8(.clk(PE_clk), .rst(rst), .in_col(sa_9_8_col), .in_row(sa_10_7_row), .out_col(sa_10_8_col), .out_row(sa_10_8_row), .out_sum(sa_out[168]));
	PE sa_10_9(.clk(PE_clk), .rst(rst), .in_col(sa_9_9_col), .in_row(sa_10_8_row), .out_col(sa_10_9_col), .out_row(sa_10_9_row), .out_sum(sa_out[169]));
	PE sa_10_10(.clk(PE_clk), .rst(rst), .in_col(sa_9_10_col), .in_row(sa_10_9_row), .out_col(sa_10_10_col), .out_row(sa_10_10_row), .out_sum(sa_out[170]));
	PE sa_10_11(.clk(PE_clk), .rst(rst), .in_col(sa_9_11_col), .in_row(sa_10_10_row), .out_col(sa_10_11_col), .out_row(sa_10_11_row), .out_sum(sa_out[171]));
	PE sa_10_12(.clk(PE_clk), .rst(rst), .in_col(sa_9_12_col), .in_row(sa_10_11_row), .out_col(sa_10_12_col), .out_row(sa_10_12_row), .out_sum(sa_out[172]));
	PE sa_10_13(.clk(PE_clk), .rst(rst), .in_col(sa_9_13_col), .in_row(sa_10_12_row), .out_col(sa_10_13_col), .out_row(sa_10_13_row), .out_sum(sa_out[173]));
	PE sa_10_14(.clk(PE_clk), .rst(rst), .in_col(sa_9_14_col), .in_row(sa_10_13_row), .out_col(sa_10_14_col), .out_row(sa_10_14_row), .out_sum(sa_out[174]));
	PE sa_10_15(.clk(PE_clk), .rst(rst), .in_col(sa_9_15_col), .in_row(sa_10_14_row), .out_col(sa_10_15_col), .out_row(sa_10_15_row), .out_sum(sa_out[175]));
	PE sa_11_0(.clk(PE_clk), .rst(rst), .in_col(sa_10_0_col), .in_row(shifter_row_11), .out_col(sa_11_0_col), .out_row(sa_11_0_row), .out_sum(sa_out[176]));
	PE sa_11_1(.clk(PE_clk), .rst(rst), .in_col(sa_10_1_col), .in_row(sa_11_0_row), .out_col(sa_11_1_col), .out_row(sa_11_1_row), .out_sum(sa_out[177]));
	PE sa_11_2(.clk(PE_clk), .rst(rst), .in_col(sa_10_2_col), .in_row(sa_11_1_row), .out_col(sa_11_2_col), .out_row(sa_11_2_row), .out_sum(sa_out[178]));
	PE sa_11_3(.clk(PE_clk), .rst(rst), .in_col(sa_10_3_col), .in_row(sa_11_2_row), .out_col(sa_11_3_col), .out_row(sa_11_3_row), .out_sum(sa_out[179]));
	PE sa_11_4(.clk(PE_clk), .rst(rst), .in_col(sa_10_4_col), .in_row(sa_11_3_row), .out_col(sa_11_4_col), .out_row(sa_11_4_row), .out_sum(sa_out[180]));
	PE sa_11_5(.clk(PE_clk), .rst(rst), .in_col(sa_10_5_col), .in_row(sa_11_4_row), .out_col(sa_11_5_col), .out_row(sa_11_5_row), .out_sum(sa_out[181]));
	PE sa_11_6(.clk(PE_clk), .rst(rst), .in_col(sa_10_6_col), .in_row(sa_11_5_row), .out_col(sa_11_6_col), .out_row(sa_11_6_row), .out_sum(sa_out[182]));
	PE sa_11_7(.clk(PE_clk), .rst(rst), .in_col(sa_10_7_col), .in_row(sa_11_6_row), .out_col(sa_11_7_col), .out_row(sa_11_7_row), .out_sum(sa_out[183]));
	PE sa_11_8(.clk(PE_clk), .rst(rst), .in_col(sa_10_8_col), .in_row(sa_11_7_row), .out_col(sa_11_8_col), .out_row(sa_11_8_row), .out_sum(sa_out[184]));
	PE sa_11_9(.clk(PE_clk), .rst(rst), .in_col(sa_10_9_col), .in_row(sa_11_8_row), .out_col(sa_11_9_col), .out_row(sa_11_9_row), .out_sum(sa_out[185]));
	PE sa_11_10(.clk(PE_clk), .rst(rst), .in_col(sa_10_10_col), .in_row(sa_11_9_row), .out_col(sa_11_10_col), .out_row(sa_11_10_row), .out_sum(sa_out[186]));
	PE sa_11_11(.clk(PE_clk), .rst(rst), .in_col(sa_10_11_col), .in_row(sa_11_10_row), .out_col(sa_11_11_col), .out_row(sa_11_11_row), .out_sum(sa_out[187]));
	PE sa_11_12(.clk(PE_clk), .rst(rst), .in_col(sa_10_12_col), .in_row(sa_11_11_row), .out_col(sa_11_12_col), .out_row(sa_11_12_row), .out_sum(sa_out[188]));
	PE sa_11_13(.clk(PE_clk), .rst(rst), .in_col(sa_10_13_col), .in_row(sa_11_12_row), .out_col(sa_11_13_col), .out_row(sa_11_13_row), .out_sum(sa_out[189]));
	PE sa_11_14(.clk(PE_clk), .rst(rst), .in_col(sa_10_14_col), .in_row(sa_11_13_row), .out_col(sa_11_14_col), .out_row(sa_11_14_row), .out_sum(sa_out[190]));
	PE sa_11_15(.clk(PE_clk), .rst(rst), .in_col(sa_10_15_col), .in_row(sa_11_14_row), .out_col(sa_11_15_col), .out_row(sa_11_15_row), .out_sum(sa_out[191]));
	PE sa_12_0(.clk(PE_clk), .rst(rst), .in_col(sa_11_0_col), .in_row(shifter_row_12), .out_col(sa_12_0_col), .out_row(sa_12_0_row), .out_sum(sa_out[192]));
	PE sa_12_1(.clk(PE_clk), .rst(rst), .in_col(sa_11_1_col), .in_row(sa_12_0_row), .out_col(sa_12_1_col), .out_row(sa_12_1_row), .out_sum(sa_out[193]));
	PE sa_12_2(.clk(PE_clk), .rst(rst), .in_col(sa_11_2_col), .in_row(sa_12_1_row), .out_col(sa_12_2_col), .out_row(sa_12_2_row), .out_sum(sa_out[194]));
	PE sa_12_3(.clk(PE_clk), .rst(rst), .in_col(sa_11_3_col), .in_row(sa_12_2_row), .out_col(sa_12_3_col), .out_row(sa_12_3_row), .out_sum(sa_out[195]));
	PE sa_12_4(.clk(PE_clk), .rst(rst), .in_col(sa_11_4_col), .in_row(sa_12_3_row), .out_col(sa_12_4_col), .out_row(sa_12_4_row), .out_sum(sa_out[196]));
	PE sa_12_5(.clk(PE_clk), .rst(rst), .in_col(sa_11_5_col), .in_row(sa_12_4_row), .out_col(sa_12_5_col), .out_row(sa_12_5_row), .out_sum(sa_out[197]));
	PE sa_12_6(.clk(PE_clk), .rst(rst), .in_col(sa_11_6_col), .in_row(sa_12_5_row), .out_col(sa_12_6_col), .out_row(sa_12_6_row), .out_sum(sa_out[198]));
	PE sa_12_7(.clk(PE_clk), .rst(rst), .in_col(sa_11_7_col), .in_row(sa_12_6_row), .out_col(sa_12_7_col), .out_row(sa_12_7_row), .out_sum(sa_out[199]));
	PE sa_12_8(.clk(PE_clk), .rst(rst), .in_col(sa_11_8_col), .in_row(sa_12_7_row), .out_col(sa_12_8_col), .out_row(sa_12_8_row), .out_sum(sa_out[200]));
	PE sa_12_9(.clk(PE_clk), .rst(rst), .in_col(sa_11_9_col), .in_row(sa_12_8_row), .out_col(sa_12_9_col), .out_row(sa_12_9_row), .out_sum(sa_out[201]));
	PE sa_12_10(.clk(PE_clk), .rst(rst), .in_col(sa_11_10_col), .in_row(sa_12_9_row), .out_col(sa_12_10_col), .out_row(sa_12_10_row), .out_sum(sa_out[202]));
	PE sa_12_11(.clk(PE_clk), .rst(rst), .in_col(sa_11_11_col), .in_row(sa_12_10_row), .out_col(sa_12_11_col), .out_row(sa_12_11_row), .out_sum(sa_out[203]));
	PE sa_12_12(.clk(PE_clk), .rst(rst), .in_col(sa_11_12_col), .in_row(sa_12_11_row), .out_col(sa_12_12_col), .out_row(sa_12_12_row), .out_sum(sa_out[204]));
	PE sa_12_13(.clk(PE_clk), .rst(rst), .in_col(sa_11_13_col), .in_row(sa_12_12_row), .out_col(sa_12_13_col), .out_row(sa_12_13_row), .out_sum(sa_out[205]));
	PE sa_12_14(.clk(PE_clk), .rst(rst), .in_col(sa_11_14_col), .in_row(sa_12_13_row), .out_col(sa_12_14_col), .out_row(sa_12_14_row), .out_sum(sa_out[206]));
	PE sa_12_15(.clk(PE_clk), .rst(rst), .in_col(sa_11_15_col), .in_row(sa_12_14_row), .out_col(sa_12_15_col), .out_row(sa_12_15_row), .out_sum(sa_out[207]));
	PE sa_13_0(.clk(PE_clk), .rst(rst), .in_col(sa_12_0_col), .in_row(shifter_row_13), .out_col(sa_13_0_col), .out_row(sa_13_0_row), .out_sum(sa_out[208]));
	PE sa_13_1(.clk(PE_clk), .rst(rst), .in_col(sa_12_1_col), .in_row(sa_13_0_row), .out_col(sa_13_1_col), .out_row(sa_13_1_row), .out_sum(sa_out[209]));
	PE sa_13_2(.clk(PE_clk), .rst(rst), .in_col(sa_12_2_col), .in_row(sa_13_1_row), .out_col(sa_13_2_col), .out_row(sa_13_2_row), .out_sum(sa_out[210]));
	PE sa_13_3(.clk(PE_clk), .rst(rst), .in_col(sa_12_3_col), .in_row(sa_13_2_row), .out_col(sa_13_3_col), .out_row(sa_13_3_row), .out_sum(sa_out[211]));
	PE sa_13_4(.clk(PE_clk), .rst(rst), .in_col(sa_12_4_col), .in_row(sa_13_3_row), .out_col(sa_13_4_col), .out_row(sa_13_4_row), .out_sum(sa_out[212]));
	PE sa_13_5(.clk(PE_clk), .rst(rst), .in_col(sa_12_5_col), .in_row(sa_13_4_row), .out_col(sa_13_5_col), .out_row(sa_13_5_row), .out_sum(sa_out[213]));
	PE sa_13_6(.clk(PE_clk), .rst(rst), .in_col(sa_12_6_col), .in_row(sa_13_5_row), .out_col(sa_13_6_col), .out_row(sa_13_6_row), .out_sum(sa_out[214]));
	PE sa_13_7(.clk(PE_clk), .rst(rst), .in_col(sa_12_7_col), .in_row(sa_13_6_row), .out_col(sa_13_7_col), .out_row(sa_13_7_row), .out_sum(sa_out[215]));
	PE sa_13_8(.clk(PE_clk), .rst(rst), .in_col(sa_12_8_col), .in_row(sa_13_7_row), .out_col(sa_13_8_col), .out_row(sa_13_8_row), .out_sum(sa_out[216]));
	PE sa_13_9(.clk(PE_clk), .rst(rst), .in_col(sa_12_9_col), .in_row(sa_13_8_row), .out_col(sa_13_9_col), .out_row(sa_13_9_row), .out_sum(sa_out[217]));
	PE sa_13_10(.clk(PE_clk), .rst(rst), .in_col(sa_12_10_col), .in_row(sa_13_9_row), .out_col(sa_13_10_col), .out_row(sa_13_10_row), .out_sum(sa_out[218]));
	PE sa_13_11(.clk(PE_clk), .rst(rst), .in_col(sa_12_11_col), .in_row(sa_13_10_row), .out_col(sa_13_11_col), .out_row(sa_13_11_row), .out_sum(sa_out[219]));
	PE sa_13_12(.clk(PE_clk), .rst(rst), .in_col(sa_12_12_col), .in_row(sa_13_11_row), .out_col(sa_13_12_col), .out_row(sa_13_12_row), .out_sum(sa_out[220]));
	PE sa_13_13(.clk(PE_clk), .rst(rst), .in_col(sa_12_13_col), .in_row(sa_13_12_row), .out_col(sa_13_13_col), .out_row(sa_13_13_row), .out_sum(sa_out[221]));
	PE sa_13_14(.clk(PE_clk), .rst(rst), .in_col(sa_12_14_col), .in_row(sa_13_13_row), .out_col(sa_13_14_col), .out_row(sa_13_14_row), .out_sum(sa_out[222]));
	PE sa_13_15(.clk(PE_clk), .rst(rst), .in_col(sa_12_15_col), .in_row(sa_13_14_row), .out_col(sa_13_15_col), .out_row(sa_13_15_row), .out_sum(sa_out[223]));
	PE sa_14_0(.clk(PE_clk), .rst(rst), .in_col(sa_13_0_col), .in_row(shifter_row_14), .out_col(sa_14_0_col), .out_row(sa_14_0_row), .out_sum(sa_out[224]));
	PE sa_14_1(.clk(PE_clk), .rst(rst), .in_col(sa_13_1_col), .in_row(sa_14_0_row), .out_col(sa_14_1_col), .out_row(sa_14_1_row), .out_sum(sa_out[225]));
	PE sa_14_2(.clk(PE_clk), .rst(rst), .in_col(sa_13_2_col), .in_row(sa_14_1_row), .out_col(sa_14_2_col), .out_row(sa_14_2_row), .out_sum(sa_out[226]));
	PE sa_14_3(.clk(PE_clk), .rst(rst), .in_col(sa_13_3_col), .in_row(sa_14_2_row), .out_col(sa_14_3_col), .out_row(sa_14_3_row), .out_sum(sa_out[227]));
	PE sa_14_4(.clk(PE_clk), .rst(rst), .in_col(sa_13_4_col), .in_row(sa_14_3_row), .out_col(sa_14_4_col), .out_row(sa_14_4_row), .out_sum(sa_out[228]));
	PE sa_14_5(.clk(PE_clk), .rst(rst), .in_col(sa_13_5_col), .in_row(sa_14_4_row), .out_col(sa_14_5_col), .out_row(sa_14_5_row), .out_sum(sa_out[229]));
	PE sa_14_6(.clk(PE_clk), .rst(rst), .in_col(sa_13_6_col), .in_row(sa_14_5_row), .out_col(sa_14_6_col), .out_row(sa_14_6_row), .out_sum(sa_out[230]));
	PE sa_14_7(.clk(PE_clk), .rst(rst), .in_col(sa_13_7_col), .in_row(sa_14_6_row), .out_col(sa_14_7_col), .out_row(sa_14_7_row), .out_sum(sa_out[231]));
	PE sa_14_8(.clk(PE_clk), .rst(rst), .in_col(sa_13_8_col), .in_row(sa_14_7_row), .out_col(sa_14_8_col), .out_row(sa_14_8_row), .out_sum(sa_out[232]));
	PE sa_14_9(.clk(PE_clk), .rst(rst), .in_col(sa_13_9_col), .in_row(sa_14_8_row), .out_col(sa_14_9_col), .out_row(sa_14_9_row), .out_sum(sa_out[233]));
	PE sa_14_10(.clk(PE_clk), .rst(rst), .in_col(sa_13_10_col), .in_row(sa_14_9_row), .out_col(sa_14_10_col), .out_row(sa_14_10_row), .out_sum(sa_out[234]));
	PE sa_14_11(.clk(PE_clk), .rst(rst), .in_col(sa_13_11_col), .in_row(sa_14_10_row), .out_col(sa_14_11_col), .out_row(sa_14_11_row), .out_sum(sa_out[235]));
	PE sa_14_12(.clk(PE_clk), .rst(rst), .in_col(sa_13_12_col), .in_row(sa_14_11_row), .out_col(sa_14_12_col), .out_row(sa_14_12_row), .out_sum(sa_out[236]));
	PE sa_14_13(.clk(PE_clk), .rst(rst), .in_col(sa_13_13_col), .in_row(sa_14_12_row), .out_col(sa_14_13_col), .out_row(sa_14_13_row), .out_sum(sa_out[237]));
	PE sa_14_14(.clk(PE_clk), .rst(rst), .in_col(sa_13_14_col), .in_row(sa_14_13_row), .out_col(sa_14_14_col), .out_row(sa_14_14_row), .out_sum(sa_out[238]));
	PE sa_14_15(.clk(PE_clk), .rst(rst), .in_col(sa_13_15_col), .in_row(sa_14_14_row), .out_col(sa_14_15_col), .out_row(sa_14_15_row), .out_sum(sa_out[239]));
	PE sa_15_0(.clk(PE_clk), .rst(rst), .in_col(sa_14_0_col), .in_row(shifter_row_15), .out_col(sa_15_0_col), .out_row(sa_15_0_row), .out_sum(sa_out[240]));
	PE sa_15_1(.clk(PE_clk), .rst(rst), .in_col(sa_14_1_col), .in_row(sa_15_0_row), .out_col(sa_15_1_col), .out_row(sa_15_1_row), .out_sum(sa_out[241]));
	PE sa_15_2(.clk(PE_clk), .rst(rst), .in_col(sa_14_2_col), .in_row(sa_15_1_row), .out_col(sa_15_2_col), .out_row(sa_15_2_row), .out_sum(sa_out[242]));
	PE sa_15_3(.clk(PE_clk), .rst(rst), .in_col(sa_14_3_col), .in_row(sa_15_2_row), .out_col(sa_15_3_col), .out_row(sa_15_3_row), .out_sum(sa_out[243]));
	PE sa_15_4(.clk(PE_clk), .rst(rst), .in_col(sa_14_4_col), .in_row(sa_15_3_row), .out_col(sa_15_4_col), .out_row(sa_15_4_row), .out_sum(sa_out[244]));
	PE sa_15_5(.clk(PE_clk), .rst(rst), .in_col(sa_14_5_col), .in_row(sa_15_4_row), .out_col(sa_15_5_col), .out_row(sa_15_5_row), .out_sum(sa_out[245]));
	PE sa_15_6(.clk(PE_clk), .rst(rst), .in_col(sa_14_6_col), .in_row(sa_15_5_row), .out_col(sa_15_6_col), .out_row(sa_15_6_row), .out_sum(sa_out[246]));
	PE sa_15_7(.clk(PE_clk), .rst(rst), .in_col(sa_14_7_col), .in_row(sa_15_6_row), .out_col(sa_15_7_col), .out_row(sa_15_7_row), .out_sum(sa_out[247]));
	PE sa_15_8(.clk(PE_clk), .rst(rst), .in_col(sa_14_8_col), .in_row(sa_15_7_row), .out_col(sa_15_8_col), .out_row(sa_15_8_row), .out_sum(sa_out[248]));
	PE sa_15_9(.clk(PE_clk), .rst(rst), .in_col(sa_14_9_col), .in_row(sa_15_8_row), .out_col(sa_15_9_col), .out_row(sa_15_9_row), .out_sum(sa_out[249]));
	PE sa_15_10(.clk(PE_clk), .rst(rst), .in_col(sa_14_10_col), .in_row(sa_15_9_row), .out_col(sa_15_10_col), .out_row(sa_15_10_row), .out_sum(sa_out[250]));
	PE sa_15_11(.clk(PE_clk), .rst(rst), .in_col(sa_14_11_col), .in_row(sa_15_10_row), .out_col(sa_15_11_col), .out_row(sa_15_11_row), .out_sum(sa_out[251]));
	PE sa_15_12(.clk(PE_clk), .rst(rst), .in_col(sa_14_12_col), .in_row(sa_15_11_row), .out_col(sa_15_12_col), .out_row(sa_15_12_row), .out_sum(sa_out[252]));
	PE sa_15_13(.clk(PE_clk), .rst(rst), .in_col(sa_14_13_col), .in_row(sa_15_12_row), .out_col(sa_15_13_col), .out_row(sa_15_13_row), .out_sum(sa_out[253]));
	PE sa_15_14(.clk(PE_clk), .rst(rst), .in_col(sa_14_14_col), .in_row(sa_15_13_row), .out_col(sa_15_14_col), .out_row(sa_15_14_row), .out_sum(sa_out[254]));
	PE sa_15_15(.clk(PE_clk), .rst(rst), .in_col(sa_14_15_col), .in_row(sa_15_14_row), .out_col(sa_15_15_col), .out_row(sa_15_15_row), .out_sum(sa_out[255]));

	// gen output addr
	reg out;

	reg finish;
	reg [7:0] oaddr;
	always @(posedge clk32x) begin
		if (row_shifter_en == 16'h0 && col_shifter_en == 16'h0 ) begin
			out <= 1;
		end
	end

	always @(posedge clk) begin
		if (oaddr == 8'd255) begin
			finish <= 1;
		end

		if (out) begin
			oaddr <= oaddr + 1;
		end
	end
	assign mc_en = 1;
	assign mc_we = out;
	assign mc_addr = oaddr;
	assign mc_din = sa_out[oaddr];
	assign ready = finish;

endmodule
